`timescale 1ns/1ps

module toplevel ( input a, output b);
    assign a = b;
endmodule

